module calculator(input wire [7:0] number, output wire [7:0] result);
    assign result = number * 2;
endmodule
